`define USE_STRUCTURAL_IMPLEMENTATION
